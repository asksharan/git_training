Hi. Welcome to the world of Mac
